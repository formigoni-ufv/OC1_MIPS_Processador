module instructionMemory (
  address,
  instruction
);

  input      [31:0] address;
  output reg [31:0] instruction;

  reg[31:0] memory[0:300];

  /*
  add $t0, $s1, $s2
  sub $t1, $s3, $s4
  beq $s5, $s6, pular
  or $s5, $t0, $t1
  slt $t3, $s1, $s2
  and $t4, $s2, $s1
  sw $t4, 4($s0)
  lw $t5, 4($s0)
  add $t6, $t4, $t5
  beq $s7, $s6, pular
  add $t0, $s1, $s2
  sub $t1, $s3, $s4
  or $s5, $t0, $t1
  slt $t3, $s1, $s2
  and $t4, $s2, $s1
  sw $t4, 0($s0)
  lw $t5, 0($s0)
  add $t6, $t4, $t5
  pular:
  add $t4, $zero, $s1
  sw $t4, 8($s0)
  lw $t5, 8($s0)
  add $t6, $t5, $t4
  */

  initial begin
        memory[ 0] = 32'b00000010001100100100000000100000;
        memory[ 4] = 32'b00000010011101000100100000100010;
        memory[ 8] = 32'b00010010101101100000000000001111;
        memory[12] = 32'b00000001000010011010100000100101;
        memory[16] = 32'b00000010001100100101100000101010;
        memory[20] = 32'b00000010010100010110000000100100;
        memory[24] = 32'b10101110000011000000000000000100;
        memory[28] = 32'b10001110000011010000000000000100;
        memory[32] = 32'b00000001100011010111000000100000;
        memory[36] = 32'b00010010111101100000000000001000;//
        memory[40] = 32'b00000010001100100100000000100000;
        memory[44] = 32'b00000010011101000100100000100010;
        memory[48] = 32'b00000001000010011010100000100101;
        memory[52] = 32'b00000010001100100101100000101010;
        memory[56] = 32'b00000010010100010110000000100100;
        memory[60] = 32'b10101110000011000000000000000000;
        memory[64] = 32'b10001110000011010000000000000000;
        memory[68] = 32'b00000001100011010111000000100000;
        memory[72] = 32'b00000000000100010110000000100000;//
        memory[76] = 32'b10101110000011000000000000001000;
        memory[80] = 32'b10001110000011010000000000001000;
        memory[84] = 32'b00000001101011000111000000100000;
    end

  always @ (address) begin
    instruction = memory[address];
  end

endmodule // instructionMemory
